module CSA_8(a1,b1,cin,sum,cout);
	input [7:0] a1,b1;
	input cin;
	output [7:0] sum;
	output cout;
	
	wire [3:0] s0,s1;
	wire c0,c1;
	wire cs;
	
	//RCA(A,B,cin,s,cout);
	RCA RCA_1(a1[3:0],b1[3:0],cin,sum[3:0],cs);
	RCA RCA_2(a1[7:4],b1[7:4],1'b0,s0[3:0],c0);
	RCA RCA_3(a1[7:4],b1[7:4],1'b1,s1[3:0],c1);
	
	//MUX
	MUX4 MUX4_1(sum[7:4],s1[3:0],s0[3:0],cs);
	//mux mux_1(cout,cs,c1,c0);
	mux mux_1(c0,c1,cs,cout);
	

endmodule

